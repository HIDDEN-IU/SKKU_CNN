`timescale 1ns/1ns
module UNPOOLING_tb();

reg CLK, RESET_N, UNPOOL_START;
reg signed [15:0] POOLED_VALUE;
reg signed [2:0] HISTORY_VALUE;

wire [15:0] UNPOOLED_VALUE;
wire UNPOOL_END, OUT_END;


initial
begin
CLK = 0;
end

initial
begin
	forever
	begin
		#5 CLK = !CLK;
	end
end

UNPOOLING #(
.SIZE(4'd8)) unpooling(
.clk(CLK),
.reset_n(RESET_N),
.unpool_start(UNPOOL_START),
.history_value(HISTORY_VALUE),
.pooled_value(POOLED_VALUE),

.unpooled_value(UNPOOLED_VALUE),
.unpool_end(UNPOOL_END),
.out_end(OUT_END)
);

initial
begin
	RESET_N = 1'b0; UNPOOL_START = 1'b0;
	#10 RESET_N = 1'b1;
    #10 UNPOOL_START = 1'b1;
    #15 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd200;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd712;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd768;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd768;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd506;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd50;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd200;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd506;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd593;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd544;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd719;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd256;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd327;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd248;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd320;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd527;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd209;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd456;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd712;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd649;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd202;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd257;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd120;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd377;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd2;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd73;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd208;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd456;
    #10 HISTORY_VALUE = 2'd2; POOLED_VALUE = 15'd712;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd338;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd3; POOLED_VALUE = 15'd376;
    #10 HISTORY_VALUE = 2'd1; POOLED_VALUE = 15'd712;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd513;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd50;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    #10 HISTORY_VALUE = 2'd0; POOLED_VALUE = 15'd0;
    
    #5000;
    $stop;
end
endmodule