module CONV_TOP(
);

endmodule