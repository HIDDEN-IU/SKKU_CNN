`timescale 1ns/1ns
module TOP_MODULE_FC_tb_R();

parameter FRT_CELL = 32;
parameter MID_CELL = 20;
parameter BCK_CELL = 10;

reg CLK, RESET_N, ENABLE, BCK_PROP_START;
reg WE, WEIGHT1, WEIGHT2, RIGHT_ANSWER, BATCH_END;
reg [15:0] ex_value, ex_addr;

wire ALL_END, FC_BCK_PROP_END, FC_BATCH_END;
wire [15:0] FC_ERR_PROP, FC_ERR_ADDR;

integer signed i, j;

initial
begin
CLK = 0;
end

initial
begin
	forever
	begin
		#5 CLK = !CLK;
	end
end

TOP_MODULE_FC #(
.FRT_CELL(FRT_CELL),
.MID_CELL(MID_CELL),
.BCK_CELL(BCK_CELL)) FC_PART(
.clk(CLK),
.reset_n(RESET_N),
.enable(ENABLE),                    //FC start when 1
.ex_we(WE),                         //flatten input write enable
.ex_value(ex_value),                //flatten input data
.ex_addr(ex_addr),                  //flatten input address
.bck_prop_start(BCK_PROP_START),    //back propagation start when 1
.batch_end(BATCH_END),              //32 mini batch finished
.weight1(WEIGHT1),                  //FC weight1 in when 1
.weight2(WEIGHT2),                  //FC weight2 in when 1
.right_answer(RIGHT_ANSWER),        //final 10 right answer when 1

.all_end(ALL_END),                  //signal to controller, FC finished when 1
.fc_bck_prop_end(FC_BCK_PROP_END),  //propagation in FC finished when 1
.fc_err_prop(FC_ERR_PROP),          //propagation error from final result
.fc_err_addr(FC_ERR_ADDR),           //propagation address
.fc_batch_end(FC_BATCH_END)
);

initial
begin
	RESET_N = 1'b0; ENABLE = 1'b0; BCK_PROP_START = 1'b0;
	#10 RESET_N = 1'b1;
    //input flatten value at ram0
    #10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b0;
    WE = 1'b1;
    #10 ex_value = 7278; ex_addr = 0;
    #10 ex_value = 5262; ex_addr = 1;
    #10 ex_value = 114; ex_addr = 2;
    #10 ex_value = 6307; ex_addr = 3;
    #10 ex_value = 74; ex_addr = 4;
    #10 ex_value = 475; ex_addr = 5;
    #10 ex_value = 2825; ex_addr = 6;
    #10 ex_value = 5284; ex_addr = 7;
    #10 ex_value = 7305; ex_addr = 8;
    #10 ex_value = 2571; ex_addr = 9;
    #10 ex_value = 0; ex_addr = 10;
    #10 ex_value = 700; ex_addr = 11;
    #10 ex_value = 1278; ex_addr = 12;
    #10 ex_value = 4991; ex_addr = 13;
    #10 ex_value = 1624; ex_addr = 14;
    #10 ex_value = 268; ex_addr = 15;
    #10 ex_value = 0; ex_addr = 16;
    #10 ex_value = 10266; ex_addr = 17;
    #10 ex_value = 453; ex_addr = 18;
    #10 ex_value = 221; ex_addr = 19;
    #10 ex_value = 6578; ex_addr = 20;
    #10 ex_value = 0; ex_addr = 21;
    #10 ex_value = 54; ex_addr = 22;
    #10 ex_value = 2715; ex_addr = 23;
    #10 ex_value = 166; ex_addr = 24;
    #10 ex_value = 90; ex_addr = 25;
    #10 ex_value = 4590; ex_addr = 26;
    #10 ex_value = 247; ex_addr = 27;
    #10 ex_value = 2324; ex_addr = 28;
    #10 ex_value = 687; ex_addr = 29;
    #10 ex_value = 404; ex_addr = 30;
    #10 ex_value = 8; ex_addr = 31;
    #10 WE = 1'b0;
    
    //input weight1 at ram0
    #10 WEIGHT1 = 1'b1; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b0;
    WE = 1'b1;
    #10 ex_value = -217; ex_addr = 32;
    #10 ex_value = -63; ex_addr = 33;
    #10 ex_value = 66; ex_addr = 34;
    #10 ex_value = -8; ex_addr = 35;
    #10 ex_value = -112; ex_addr = 36;
    #10 ex_value = 249; ex_addr = 37;
    #10 ex_value = -98; ex_addr = 38;
    #10 ex_value = 200; ex_addr = 39;
    #10 ex_value = -157; ex_addr = 40;
    #10 ex_value = -52; ex_addr = 41;
    #10 ex_value = 114; ex_addr = 42;
    #10 ex_value = -8; ex_addr = 43;
    #10 ex_value = -192; ex_addr = 44;
    #10 ex_value = -203; ex_addr = 45;
    #10 ex_value = -208; ex_addr = 46;
    #10 ex_value = -190; ex_addr = 47;
    #10 ex_value = -17; ex_addr = 48;
    #10 ex_value = -147; ex_addr = 49;
    #10 ex_value = 116; ex_addr = 50;
    #10 ex_value = 110; ex_addr = 51;
    #10 ex_value = 150; ex_addr = 52;
    #10 ex_value = -138; ex_addr = 53;
    #10 ex_value = -162; ex_addr = 54;
    #10 ex_value = -28; ex_addr = 55;
    #10 ex_value = -191; ex_addr = 56;
    #10 ex_value = -45; ex_addr = 57;
    #10 ex_value = 86; ex_addr = 58;
    #10 ex_value = -110; ex_addr = 59;
    #10 ex_value = 129; ex_addr = 60;
    #10 ex_value = -142; ex_addr = 61;
    #10 ex_value = -193; ex_addr = 62;
    #10 ex_value = -4; ex_addr = 63;
    #10 ex_value = -226; ex_addr = 64;
    #10 ex_value = -143; ex_addr = 65;
    #10 ex_value = -158; ex_addr = 66;
    #10 ex_value = -117; ex_addr = 67;
    #10 ex_value = -39; ex_addr = 68;
    #10 ex_value = 205; ex_addr = 69;
    #10 ex_value = -198; ex_addr = 70;
    #10 ex_value = 214; ex_addr = 71;
    #10 ex_value = -58; ex_addr = 72;
    #10 ex_value = -160; ex_addr = 73;
    #10 ex_value = -102; ex_addr = 74;
    #10 ex_value = 38; ex_addr = 75;
    #10 ex_value = -5; ex_addr = 76;
    #10 ex_value = -158; ex_addr = 77;
    #10 ex_value = 25; ex_addr = 78;
    #10 ex_value = 2; ex_addr = 79;
    #10 ex_value = 52; ex_addr = 80;
    #10 ex_value = -145; ex_addr = 81;
    #10 ex_value = 70; ex_addr = 82;
    #10 ex_value = 0; ex_addr = 83;
    #10 ex_value = 170; ex_addr = 84;
    #10 ex_value = -45; ex_addr = 85;
    #10 ex_value = 113; ex_addr = 86;
    #10 ex_value = 171; ex_addr = 87;
    #10 ex_value = 6; ex_addr = 88;
    #10 ex_value = -19; ex_addr = 89;
    #10 ex_value = -181; ex_addr = 90;
    #10 ex_value = 29; ex_addr = 91;
    #10 ex_value = -104; ex_addr = 92;
    #10 ex_value = 97; ex_addr = 93;
    #10 ex_value = 114; ex_addr = 94;
    #10 ex_value = 83; ex_addr = 95;
    #10 ex_value = -28; ex_addr = 96;
    #10 ex_value = -119; ex_addr = 97;
    #10 ex_value = -241; ex_addr = 98;
    #10 ex_value = 119; ex_addr = 99;
    #10 ex_value = -31; ex_addr = 100;
    #10 ex_value = -7; ex_addr = 101;
    #10 ex_value = 70; ex_addr = 102;
    #10 ex_value = 6; ex_addr = 103;
    #10 ex_value = 229; ex_addr = 104;
    #10 ex_value = 238; ex_addr = 105;
    #10 ex_value = 108; ex_addr = 106;
    #10 ex_value = 30; ex_addr = 107;
    #10 ex_value = 255; ex_addr = 108;
    #10 ex_value = 35; ex_addr = 109;
    #10 ex_value = -69; ex_addr = 110;
    #10 ex_value = 133; ex_addr = 111;
    #10 ex_value = -75; ex_addr = 112;
    #10 ex_value = 88; ex_addr = 113;
    #10 ex_value = 175; ex_addr = 114;
    #10 ex_value = 121; ex_addr = 115;
    #10 ex_value = 88; ex_addr = 116;
    #10 ex_value = 57; ex_addr = 117;
    #10 ex_value = -146; ex_addr = 118;
    #10 ex_value = 31; ex_addr = 119;
    #10 ex_value = 139; ex_addr = 120;
    #10 ex_value = -172; ex_addr = 121;
    #10 ex_value = -153; ex_addr = 122;
    #10 ex_value = -165; ex_addr = 123;
    #10 ex_value = 83; ex_addr = 124;
    #10 ex_value = -204; ex_addr = 125;
    #10 ex_value = -231; ex_addr = 126;
    #10 ex_value = 173; ex_addr = 127;
    #10 ex_value = -222; ex_addr = 128;
    #10 ex_value = 97; ex_addr = 129;
    #10 ex_value = 50; ex_addr = 130;
    #10 ex_value = 248; ex_addr = 131;
    #10 ex_value = 140; ex_addr = 132;
    #10 ex_value = -80; ex_addr = 133;
    #10 ex_value = -77; ex_addr = 134;
    #10 ex_value = -181; ex_addr = 135;
    #10 ex_value = 160; ex_addr = 136;
    #10 ex_value = 52; ex_addr = 137;
    #10 ex_value = 45; ex_addr = 138;
    #10 ex_value = 15; ex_addr = 139;
    #10 ex_value = 21; ex_addr = 140;
    #10 ex_value = -246; ex_addr = 141;
    #10 ex_value = -103; ex_addr = 142;
    #10 ex_value = 154; ex_addr = 143;
    #10 ex_value = 104; ex_addr = 144;
    #10 ex_value = -101; ex_addr = 145;
    #10 ex_value = -60; ex_addr = 146;
    #10 ex_value = -14; ex_addr = 147;
    #10 ex_value = 136; ex_addr = 148;
    #10 ex_value = 61; ex_addr = 149;
    #10 ex_value = -60; ex_addr = 150;
    #10 ex_value = -104; ex_addr = 151;
    #10 ex_value = 153; ex_addr = 152;
    #10 ex_value = -156; ex_addr = 153;
    #10 ex_value = -179; ex_addr = 154;
    #10 ex_value = 67; ex_addr = 155;
    #10 ex_value = -84; ex_addr = 156;
    #10 ex_value = 191; ex_addr = 157;
    #10 ex_value = 130; ex_addr = 158;
    #10 ex_value = -33; ex_addr = 159;
    #10 ex_value = 71; ex_addr = 160;
    #10 ex_value = -151; ex_addr = 161;
    #10 ex_value = -108; ex_addr = 162;
    #10 ex_value = 143; ex_addr = 163;
    #10 ex_value = 13; ex_addr = 164;
    #10 ex_value = -46; ex_addr = 165;
    #10 ex_value = 157; ex_addr = 166;
    #10 ex_value = 244; ex_addr = 167;
    #10 ex_value = 78; ex_addr = 168;
    #10 ex_value = 189; ex_addr = 169;
    #10 ex_value = 45; ex_addr = 170;
    #10 ex_value = 154; ex_addr = 171;
    #10 ex_value = -190; ex_addr = 172;
    #10 ex_value = -228; ex_addr = 173;
    #10 ex_value = 168; ex_addr = 174;
    #10 ex_value = -90; ex_addr = 175;
    #10 ex_value = -175; ex_addr = 176;
    #10 ex_value = -10; ex_addr = 177;
    #10 ex_value = 78; ex_addr = 178;
    #10 ex_value = -81; ex_addr = 179;
    #10 ex_value = 217; ex_addr = 180;
    #10 ex_value = -107; ex_addr = 181;
    #10 ex_value = -90; ex_addr = 182;
    #10 ex_value = 120; ex_addr = 183;
    #10 ex_value = 165; ex_addr = 184;
    #10 ex_value = -167; ex_addr = 185;
    #10 ex_value = -46; ex_addr = 186;
    #10 ex_value = -55; ex_addr = 187;
    #10 ex_value = -231; ex_addr = 188;
    #10 ex_value = -28; ex_addr = 189;
    #10 ex_value = -46; ex_addr = 190;
    #10 ex_value = -59; ex_addr = 191;
    #10 ex_value = -70; ex_addr = 192;
    #10 ex_value = 154; ex_addr = 193;
    #10 ex_value = 166; ex_addr = 194;
    #10 ex_value = -53; ex_addr = 195;
    #10 ex_value = -217; ex_addr = 196;
    #10 ex_value = 242; ex_addr = 197;
    #10 ex_value = -246; ex_addr = 198;
    #10 ex_value = 213; ex_addr = 199;
    #10 ex_value = 242; ex_addr = 200;
    #10 ex_value = -53; ex_addr = 201;
    #10 ex_value = 248; ex_addr = 202;
    #10 ex_value = 110; ex_addr = 203;
    #10 ex_value = -195; ex_addr = 204;
    #10 ex_value = -128; ex_addr = 205;
    #10 ex_value = -45; ex_addr = 206;
    #10 ex_value = -255; ex_addr = 207;
    #10 ex_value = -115; ex_addr = 208;
    #10 ex_value = 99; ex_addr = 209;
    #10 ex_value = 90; ex_addr = 210;
    #10 ex_value = -171; ex_addr = 211;
    #10 ex_value = 186; ex_addr = 212;
    #10 ex_value = -195; ex_addr = 213;
    #10 ex_value = 133; ex_addr = 214;
    #10 ex_value = 128; ex_addr = 215;
    #10 ex_value = 247; ex_addr = 216;
    #10 ex_value = -189; ex_addr = 217;
    #10 ex_value = -104; ex_addr = 218;
    #10 ex_value = 225; ex_addr = 219;
    #10 ex_value = -22; ex_addr = 220;
    #10 ex_value = -107; ex_addr = 221;
    #10 ex_value = 173; ex_addr = 222;
    #10 ex_value = 82; ex_addr = 223;
    #10 ex_value = -104; ex_addr = 224;
    #10 ex_value = -12; ex_addr = 225;
    #10 ex_value = -207; ex_addr = 226;
    #10 ex_value = -193; ex_addr = 227;
    #10 ex_value = -189; ex_addr = 228;
    #10 ex_value = -45; ex_addr = 229;
    #10 ex_value = -38; ex_addr = 230;
    #10 ex_value = 167; ex_addr = 231;
    #10 ex_value = -70; ex_addr = 232;
    #10 ex_value = 157; ex_addr = 233;
    #10 ex_value = 221; ex_addr = 234;
    #10 ex_value = 138; ex_addr = 235;
    #10 ex_value = 19; ex_addr = 236;
    #10 ex_value = 105; ex_addr = 237;
    #10 ex_value = 226; ex_addr = 238;
    #10 ex_value = 136; ex_addr = 239;
    #10 ex_value = 167; ex_addr = 240;
    #10 ex_value = -59; ex_addr = 241;
    #10 ex_value = 121; ex_addr = 242;
    #10 ex_value = 252; ex_addr = 243;
    #10 ex_value = -106; ex_addr = 244;
    #10 ex_value = 117; ex_addr = 245;
    #10 ex_value = 220; ex_addr = 246;
    #10 ex_value = 112; ex_addr = 247;
    #10 ex_value = -199; ex_addr = 248;
    #10 ex_value = 140; ex_addr = 249;
    #10 ex_value = -84; ex_addr = 250;
    #10 ex_value = -58; ex_addr = 251;
    #10 ex_value = -54; ex_addr = 252;
    #10 ex_value = 77; ex_addr = 253;
    #10 ex_value = 123; ex_addr = 254;
    #10 ex_value = 199; ex_addr = 255;
    #10 ex_value = 129; ex_addr = 256;
    #10 ex_value = -107; ex_addr = 257;
    #10 ex_value = 107; ex_addr = 258;
    #10 ex_value = -84; ex_addr = 259;
    #10 ex_value = -24; ex_addr = 260;
    #10 ex_value = -30; ex_addr = 261;
    #10 ex_value = -17; ex_addr = 262;
    #10 ex_value = 122; ex_addr = 263;
    #10 ex_value = 244; ex_addr = 264;
    #10 ex_value = -250; ex_addr = 265;
    #10 ex_value = 125; ex_addr = 266;
    #10 ex_value = 111; ex_addr = 267;
    #10 ex_value = -139; ex_addr = 268;
    #10 ex_value = -188; ex_addr = 269;
    #10 ex_value = 85; ex_addr = 270;
    #10 ex_value = 249; ex_addr = 271;
    #10 ex_value = 163; ex_addr = 272;
    #10 ex_value = 210; ex_addr = 273;
    #10 ex_value = 255; ex_addr = 274;
    #10 ex_value = -10; ex_addr = 275;
    #10 ex_value = -162; ex_addr = 276;
    #10 ex_value = -188; ex_addr = 277;
    #10 ex_value = -72; ex_addr = 278;
    #10 ex_value = -57; ex_addr = 279;
    #10 ex_value = 191; ex_addr = 280;
    #10 ex_value = 139; ex_addr = 281;
    #10 ex_value = 228; ex_addr = 282;
    #10 ex_value = 18; ex_addr = 283;
    #10 ex_value = -220; ex_addr = 284;
    #10 ex_value = 84; ex_addr = 285;
    #10 ex_value = 156; ex_addr = 286;
    #10 ex_value = -55; ex_addr = 287;
    #10 ex_value = -201; ex_addr = 288;
    #10 ex_value = 60; ex_addr = 289;
    #10 ex_value = -107; ex_addr = 290;
    #10 ex_value = -215; ex_addr = 291;
    #10 ex_value = -245; ex_addr = 292;
    #10 ex_value = 136; ex_addr = 293;
    #10 ex_value = 113; ex_addr = 294;
    #10 ex_value = 44; ex_addr = 295;
    #10 ex_value = -192; ex_addr = 296;
    #10 ex_value = -245; ex_addr = 297;
    #10 ex_value = -187; ex_addr = 298;
    #10 ex_value = -96; ex_addr = 299;
    #10 ex_value = -46; ex_addr = 300;
    #10 ex_value = -137; ex_addr = 301;
    #10 ex_value = 11; ex_addr = 302;
    #10 ex_value = 55; ex_addr = 303;
    #10 ex_value = 46; ex_addr = 304;
    #10 ex_value = -122; ex_addr = 305;
    #10 ex_value = -109; ex_addr = 306;
    #10 ex_value = 7; ex_addr = 307;
    #10 ex_value = 255; ex_addr = 308;
    #10 ex_value = 75; ex_addr = 309;
    #10 ex_value = -227; ex_addr = 310;
    #10 ex_value = 203; ex_addr = 311;
    #10 ex_value = 136; ex_addr = 312;
    #10 ex_value = 172; ex_addr = 313;
    #10 ex_value = 162; ex_addr = 314;
    #10 ex_value = -230; ex_addr = 315;
    #10 ex_value = 218; ex_addr = 316;
    #10 ex_value = -227; ex_addr = 317;
    #10 ex_value = -118; ex_addr = 318;
    #10 ex_value = 189; ex_addr = 319;
    #10 ex_value = 138; ex_addr = 320;
    #10 ex_value = 67; ex_addr = 321;
    #10 ex_value = 89; ex_addr = 322;
    #10 ex_value = 15; ex_addr = 323;
    #10 ex_value = -13; ex_addr = 324;
    #10 ex_value = -111; ex_addr = 325;
    #10 ex_value = -213; ex_addr = 326;
    #10 ex_value = 36; ex_addr = 327;
    #10 ex_value = 109; ex_addr = 328;
    #10 ex_value = -160; ex_addr = 329;
    #10 ex_value = 161; ex_addr = 330;
    #10 ex_value = -226; ex_addr = 331;
    #10 ex_value = -205; ex_addr = 332;
    #10 ex_value = -238; ex_addr = 333;
    #10 ex_value = 70; ex_addr = 334;
    #10 ex_value = 45; ex_addr = 335;
    #10 ex_value = 130; ex_addr = 336;
    #10 ex_value = -133; ex_addr = 337;
    #10 ex_value = 46; ex_addr = 338;
    #10 ex_value = 88; ex_addr = 339;
    #10 ex_value = -6; ex_addr = 340;
    #10 ex_value = -80; ex_addr = 341;
    #10 ex_value = -77; ex_addr = 342;
    #10 ex_value = -80; ex_addr = 343;
    #10 ex_value = 41; ex_addr = 344;
    #10 ex_value = -189; ex_addr = 345;
    #10 ex_value = 98; ex_addr = 346;
    #10 ex_value = -215; ex_addr = 347;
    #10 ex_value = 51; ex_addr = 348;
    #10 ex_value = 129; ex_addr = 349;
    #10 ex_value = 115; ex_addr = 350;
    #10 ex_value = -40; ex_addr = 351;
    #10 ex_value = -163; ex_addr = 352;
    #10 ex_value = -106; ex_addr = 353;
    #10 ex_value = 84; ex_addr = 354;
    #10 ex_value = -158; ex_addr = 355;
    #10 ex_value = 214; ex_addr = 356;
    #10 ex_value = 48; ex_addr = 357;
    #10 ex_value = -64; ex_addr = 358;
    #10 ex_value = -42; ex_addr = 359;
    #10 ex_value = -208; ex_addr = 360;
    #10 ex_value = -182; ex_addr = 361;
    #10 ex_value = -18; ex_addr = 362;
    #10 ex_value = -182; ex_addr = 363;
    #10 ex_value = -48; ex_addr = 364;
    #10 ex_value = -33; ex_addr = 365;
    #10 ex_value = -215; ex_addr = 366;
    #10 ex_value = -235; ex_addr = 367;
    #10 ex_value = -226; ex_addr = 368;
    #10 ex_value = 88; ex_addr = 369;
    #10 ex_value = -207; ex_addr = 370;
    #10 ex_value = 6; ex_addr = 371;
    #10 ex_value = -235; ex_addr = 372;
    #10 ex_value = -118; ex_addr = 373;
    #10 ex_value = -141; ex_addr = 374;
    #10 ex_value = 84; ex_addr = 375;
    #10 ex_value = 127; ex_addr = 376;
    #10 ex_value = -7; ex_addr = 377;
    #10 ex_value = 31; ex_addr = 378;
    #10 ex_value = -229; ex_addr = 379;
    #10 ex_value = -16; ex_addr = 380;
    #10 ex_value = 25; ex_addr = 381;
    #10 ex_value = -249; ex_addr = 382;
    #10 ex_value = 183; ex_addr = 383;
    #10 ex_value = -13; ex_addr = 384;
    #10 ex_value = 239; ex_addr = 385;
    #10 ex_value = 235; ex_addr = 386;
    #10 ex_value = 198; ex_addr = 387;
    #10 ex_value = -174; ex_addr = 388;
    #10 ex_value = 142; ex_addr = 389;
    #10 ex_value = -255; ex_addr = 390;
    #10 ex_value = 206; ex_addr = 391;
    #10 ex_value = 40; ex_addr = 392;
    #10 ex_value = -176; ex_addr = 393;
    #10 ex_value = 236; ex_addr = 394;
    #10 ex_value = 37; ex_addr = 395;
    #10 ex_value = -121; ex_addr = 396;
    #10 ex_value = -190; ex_addr = 397;
    #10 ex_value = -255; ex_addr = 398;
    #10 ex_value = 155; ex_addr = 399;
    #10 ex_value = 37; ex_addr = 400;
    #10 ex_value = 205; ex_addr = 401;
    #10 ex_value = -99; ex_addr = 402;
    #10 ex_value = -237; ex_addr = 403;
    #10 ex_value = -51; ex_addr = 404;
    #10 ex_value = -53; ex_addr = 405;
    #10 ex_value = 245; ex_addr = 406;
    #10 ex_value = 142; ex_addr = 407;
    #10 ex_value = -39; ex_addr = 408;
    #10 ex_value = 206; ex_addr = 409;
    #10 ex_value = -155; ex_addr = 410;
    #10 ex_value = -66; ex_addr = 411;
    #10 ex_value = -13; ex_addr = 412;
    #10 ex_value = 156; ex_addr = 413;
    #10 ex_value = -36; ex_addr = 414;
    #10 ex_value = -6; ex_addr = 415;
    #10 ex_value = -140; ex_addr = 416;
    #10 ex_value = 254; ex_addr = 417;
    #10 ex_value = -212; ex_addr = 418;
    #10 ex_value = 234; ex_addr = 419;
    #10 ex_value = 86; ex_addr = 420;
    #10 ex_value = -27; ex_addr = 421;
    #10 ex_value = -120; ex_addr = 422;
    #10 ex_value = -11; ex_addr = 423;
    #10 ex_value = -135; ex_addr = 424;
    #10 ex_value = 119; ex_addr = 425;
    #10 ex_value = -42; ex_addr = 426;
    #10 ex_value = 173; ex_addr = 427;
    #10 ex_value = -245; ex_addr = 428;
    #10 ex_value = 255; ex_addr = 429;
    #10 ex_value = 169; ex_addr = 430;
    #10 ex_value = 37; ex_addr = 431;
    #10 ex_value = -102; ex_addr = 432;
    #10 ex_value = 173; ex_addr = 433;
    #10 ex_value = 112; ex_addr = 434;
    #10 ex_value = 110; ex_addr = 435;
    #10 ex_value = -198; ex_addr = 436;
    #10 ex_value = 173; ex_addr = 437;
    #10 ex_value = 209; ex_addr = 438;
    #10 ex_value = -227; ex_addr = 439;
    #10 ex_value = 206; ex_addr = 440;
    #10 ex_value = -202; ex_addr = 441;
    #10 ex_value = 218; ex_addr = 442;
    #10 ex_value = 13; ex_addr = 443;
    #10 ex_value = -112; ex_addr = 444;
    #10 ex_value = 222; ex_addr = 445;
    #10 ex_value = 202; ex_addr = 446;
    #10 ex_value = 75; ex_addr = 447;
    #10 ex_value = -163; ex_addr = 448;
    #10 ex_value = -239; ex_addr = 449;
    #10 ex_value = -91; ex_addr = 450;
    #10 ex_value = -238; ex_addr = 451;
    #10 ex_value = -96; ex_addr = 452;
    #10 ex_value = -125; ex_addr = 453;
    #10 ex_value = -61; ex_addr = 454;
    #10 ex_value = 50; ex_addr = 455;
    #10 ex_value = -28; ex_addr = 456;
    #10 ex_value = -181; ex_addr = 457;
    #10 ex_value = -187; ex_addr = 458;
    #10 ex_value = 72; ex_addr = 459;
    #10 ex_value = 184; ex_addr = 460;
    #10 ex_value = -66; ex_addr = 461;
    #10 ex_value = 230; ex_addr = 462;
    #10 ex_value = 161; ex_addr = 463;
    #10 ex_value = -103; ex_addr = 464;
    #10 ex_value = -141; ex_addr = 465;
    #10 ex_value = 250; ex_addr = 466;
    #10 ex_value = 216; ex_addr = 467;
    #10 ex_value = 80; ex_addr = 468;
    #10 ex_value = -249; ex_addr = 469;
    #10 ex_value = -94; ex_addr = 470;
    #10 ex_value = -93; ex_addr = 471;
    #10 ex_value = 160; ex_addr = 472;
    #10 ex_value = 38; ex_addr = 473;
    #10 ex_value = -77; ex_addr = 474;
    #10 ex_value = -156; ex_addr = 475;
    #10 ex_value = 167; ex_addr = 476;
    #10 ex_value = -181; ex_addr = 477;
    #10 ex_value = 168; ex_addr = 478;
    #10 ex_value = 77; ex_addr = 479;
    #10 ex_value = 191; ex_addr = 480;
    #10 ex_value = -9; ex_addr = 481;
    #10 ex_value = 148; ex_addr = 482;
    #10 ex_value = -123; ex_addr = 483;
    #10 ex_value = 10; ex_addr = 484;
    #10 ex_value = 137; ex_addr = 485;
    #10 ex_value = 213; ex_addr = 486;
    #10 ex_value = 127; ex_addr = 487;
    #10 ex_value = -233; ex_addr = 488;
    #10 ex_value = 152; ex_addr = 489;
    #10 ex_value = 172; ex_addr = 490;
    #10 ex_value = -16; ex_addr = 491;
    #10 ex_value = 153; ex_addr = 492;
    #10 ex_value = 231; ex_addr = 493;
    #10 ex_value = 27; ex_addr = 494;
    #10 ex_value = 155; ex_addr = 495;
    #10 ex_value = -13; ex_addr = 496;
    #10 ex_value = -173; ex_addr = 497;
    #10 ex_value = 94; ex_addr = 498;
    #10 ex_value = -93; ex_addr = 499;
    #10 ex_value = 61; ex_addr = 500;
    #10 ex_value = -239; ex_addr = 501;
    #10 ex_value = 237; ex_addr = 502;
    #10 ex_value = 119; ex_addr = 503;
    #10 ex_value = 239; ex_addr = 504;
    #10 ex_value = -41; ex_addr = 505;
    #10 ex_value = 213; ex_addr = 506;
    #10 ex_value = -74; ex_addr = 507;
    #10 ex_value = 56; ex_addr = 508;
    #10 ex_value = 111; ex_addr = 509;
    #10 ex_value = -14; ex_addr = 510;
    #10 ex_value = -152; ex_addr = 511;
    #10 ex_value = 30; ex_addr = 512;
    #10 ex_value = 169; ex_addr = 513;
    #10 ex_value = -70; ex_addr = 514;
    #10 ex_value = 168; ex_addr = 515;
    #10 ex_value = 181; ex_addr = 516;
    #10 ex_value = -92; ex_addr = 517;
    #10 ex_value = 109; ex_addr = 518;
    #10 ex_value = 138; ex_addr = 519;
    #10 ex_value = 118; ex_addr = 520;
    #10 ex_value = 4; ex_addr = 521;
    #10 ex_value = -20; ex_addr = 522;
    #10 ex_value = -240; ex_addr = 523;
    #10 ex_value = -64; ex_addr = 524;
    #10 ex_value = -198; ex_addr = 525;
    #10 ex_value = 219; ex_addr = 526;
    #10 ex_value = -117; ex_addr = 527;
    #10 ex_value = -4; ex_addr = 528;
    #10 ex_value = -10; ex_addr = 529;
    #10 ex_value = -229; ex_addr = 530;
    #10 ex_value = 225; ex_addr = 531;
    #10 ex_value = 180; ex_addr = 532;
    #10 ex_value = 7; ex_addr = 533;
    #10 ex_value = -118; ex_addr = 534;
    #10 ex_value = -21; ex_addr = 535;
    #10 ex_value = -179; ex_addr = 536;
    #10 ex_value = -140; ex_addr = 537;
    #10 ex_value = -201; ex_addr = 538;
    #10 ex_value = -99; ex_addr = 539;
    #10 ex_value = -35; ex_addr = 540;
    #10 ex_value = 135; ex_addr = 541;
    #10 ex_value = -37; ex_addr = 542;
    #10 ex_value = -112; ex_addr = 543;
    #10 ex_value = -251; ex_addr = 544;
    #10 ex_value = 155; ex_addr = 545;
    #10 ex_value = 163; ex_addr = 546;
    #10 ex_value = -54; ex_addr = 547;
    #10 ex_value = -60; ex_addr = 548;
    #10 ex_value = -104; ex_addr = 549;
    #10 ex_value = 179; ex_addr = 550;
    #10 ex_value = 28; ex_addr = 551;
    #10 ex_value = -8; ex_addr = 552;
    #10 ex_value = -57; ex_addr = 553;
    #10 ex_value = -57; ex_addr = 554;
    #10 ex_value = -97; ex_addr = 555;
    #10 ex_value = 89; ex_addr = 556;
    #10 ex_value = 104; ex_addr = 557;
    #10 ex_value = 195; ex_addr = 558;
    #10 ex_value = 245; ex_addr = 559;
    #10 ex_value = 203; ex_addr = 560;
    #10 ex_value = 121; ex_addr = 561;
    #10 ex_value = -218; ex_addr = 562;
    #10 ex_value = 154; ex_addr = 563;
    #10 ex_value = 255; ex_addr = 564;
    #10 ex_value = 230; ex_addr = 565;
    #10 ex_value = -61; ex_addr = 566;
    #10 ex_value = -188; ex_addr = 567;
    #10 ex_value = -224; ex_addr = 568;
    #10 ex_value = 165; ex_addr = 569;
    #10 ex_value = -223; ex_addr = 570;
    #10 ex_value = -247; ex_addr = 571;
    #10 ex_value = -104; ex_addr = 572;
    #10 ex_value = -47; ex_addr = 573;
    #10 ex_value = -125; ex_addr = 574;
    #10 ex_value = 114; ex_addr = 575;
    #10 ex_value = 95; ex_addr = 576;
    #10 ex_value = -231; ex_addr = 577;
    #10 ex_value = -126; ex_addr = 578;
    #10 ex_value = 6; ex_addr = 579;
    #10 ex_value = 117; ex_addr = 580;
    #10 ex_value = 195; ex_addr = 581;
    #10 ex_value = 74; ex_addr = 582;
    #10 ex_value = -110; ex_addr = 583;
    #10 ex_value = 58; ex_addr = 584;
    #10 ex_value = 114; ex_addr = 585;
    #10 ex_value = 156; ex_addr = 586;
    #10 ex_value = 107; ex_addr = 587;
    #10 ex_value = 99; ex_addr = 588;
    #10 ex_value = 170; ex_addr = 589;
    #10 ex_value = -201; ex_addr = 590;
    #10 ex_value = 58; ex_addr = 591;
    #10 ex_value = 203; ex_addr = 592;
    #10 ex_value = -225; ex_addr = 593;
    #10 ex_value = 255; ex_addr = 594;
    #10 ex_value = 189; ex_addr = 595;
    #10 ex_value = -188; ex_addr = 596;
    #10 ex_value = -97; ex_addr = 597;
    #10 ex_value = 243; ex_addr = 598;
    #10 ex_value = 168; ex_addr = 599;
    #10 ex_value = 245; ex_addr = 600;
    #10 ex_value = -246; ex_addr = 601;
    #10 ex_value = 102; ex_addr = 602;
    #10 ex_value = 254; ex_addr = 603;
    #10 ex_value = -83; ex_addr = 604;
    #10 ex_value = -101; ex_addr = 605;
    #10 ex_value = 74; ex_addr = 606;
    #10 ex_value = 255; ex_addr = 607;
    #10 ex_value = 242; ex_addr = 608;
    #10 ex_value = -165; ex_addr = 609;
    #10 ex_value = -160; ex_addr = 610;
    #10 ex_value = -232; ex_addr = 611;
    #10 ex_value = 178; ex_addr = 612;
    #10 ex_value = -103; ex_addr = 613;
    #10 ex_value = 115; ex_addr = 614;
    #10 ex_value = -46; ex_addr = 615;
    #10 ex_value = 63; ex_addr = 616;
    #10 ex_value = 52; ex_addr = 617;
    #10 ex_value = -253; ex_addr = 618;
    #10 ex_value = -222; ex_addr = 619;
    #10 ex_value = -36; ex_addr = 620;
    #10 ex_value = -28; ex_addr = 621;
    #10 ex_value = -45; ex_addr = 622;
    #10 ex_value = 221; ex_addr = 623;
    #10 ex_value = 240; ex_addr = 624;
    #10 ex_value = 27; ex_addr = 625;
    #10 ex_value = 234; ex_addr = 626;
    #10 ex_value = -68; ex_addr = 627;
    #10 ex_value = 172; ex_addr = 628;
    #10 ex_value = 181; ex_addr = 629;
    #10 ex_value = -100; ex_addr = 630;
    #10 ex_value = 113; ex_addr = 631;
    #10 ex_value = 124; ex_addr = 632;
    #10 ex_value = -188; ex_addr = 633;
    #10 ex_value = -233; ex_addr = 634;
    #10 ex_value = 147; ex_addr = 635;
    #10 ex_value = 18; ex_addr = 636;
    #10 ex_value = -132; ex_addr = 637;
    #10 ex_value = -116; ex_addr = 638;
    #10 ex_value = 6; ex_addr = 639;
    #10 ex_value = 29; ex_addr = 640;
    #10 ex_value = 214; ex_addr = 641;
    #10 ex_value = 233; ex_addr = 642;
    #10 ex_value = -163; ex_addr = 643;
    #10 ex_value = 220; ex_addr = 644;
    #10 ex_value = -2; ex_addr = 645;
    #10 ex_value = 13; ex_addr = 646;
    #10 ex_value = -73; ex_addr = 647;
    #10 ex_value = -25; ex_addr = 648;
    #10 ex_value = -101; ex_addr = 649;
    #10 ex_value = 206; ex_addr = 650;
    #10 ex_value = 111; ex_addr = 651;
    #10 ex_value = -97; ex_addr = 652;
    #10 ex_value = -230; ex_addr = 653;
    #10 ex_value = 122; ex_addr = 654;
    #10 ex_value = -48; ex_addr = 655;
    #10 ex_value = 169; ex_addr = 656;
    #10 ex_value = -89; ex_addr = 657;
    #10 ex_value = -197; ex_addr = 658;
    #10 ex_value = 5; ex_addr = 659;
    #10 ex_value = 114; ex_addr = 660;
    #10 ex_value = 6; ex_addr = 661;
    #10 ex_value = 100; ex_addr = 662;
    #10 ex_value = -20; ex_addr = 663;
    #10 ex_value = -54; ex_addr = 664;
    #10 ex_value = 146; ex_addr = 665;
    #10 ex_value = -169; ex_addr = 666;
    #10 ex_value = 49; ex_addr = 667;
    #10 ex_value = 158; ex_addr = 668;
    #10 ex_value = -62; ex_addr = 669;
    #10 ex_value = 175; ex_addr = 670;
    #10 ex_value = 224; ex_addr = 671;
    #10 WE = 1'b0;
    
    //input weight2 at ram1
    #10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b1; RIGHT_ANSWER = 1'b0;
    WE = 1'b1;
    #10 ex_value = 184; ex_addr = 20;
    #10 ex_value = -10; ex_addr = 21;
    #10 ex_value = 42; ex_addr = 22;
    #10 ex_value = 73; ex_addr = 23;
    #10 ex_value = -42; ex_addr = 24;
    #10 ex_value = -14; ex_addr = 25;
    #10 ex_value = 190; ex_addr = 26;
    #10 ex_value = 35; ex_addr = 27;
    #10 ex_value = -45; ex_addr = 28;
    #10 ex_value = -195; ex_addr = 29;
    #10 ex_value = 104; ex_addr = 30;
    #10 ex_value = 233; ex_addr = 31;
    #10 ex_value = 48; ex_addr = 32;
    #10 ex_value = -220; ex_addr = 33;
    #10 ex_value = -182; ex_addr = 34;
    #10 ex_value = -11; ex_addr = 35;
    #10 ex_value = -124; ex_addr = 36;
    #10 ex_value = -7; ex_addr = 37;
    #10 ex_value = -171; ex_addr = 38;
    #10 ex_value = 249; ex_addr = 39;
    #10 ex_value = -204; ex_addr = 40;
    #10 ex_value = 110; ex_addr = 41;
    #10 ex_value = -57; ex_addr = 42;
    #10 ex_value = -240; ex_addr = 43;
    #10 ex_value = -16; ex_addr = 44;
    #10 ex_value = 233; ex_addr = 45;
    #10 ex_value = -226; ex_addr = 46;
    #10 ex_value = 72; ex_addr = 47;
    #10 ex_value = 6; ex_addr = 48;
    #10 ex_value = -218; ex_addr = 49;
    #10 ex_value = 11; ex_addr = 50;
    #10 ex_value = -53; ex_addr = 51;
    #10 ex_value = -29; ex_addr = 52;
    #10 ex_value = -217; ex_addr = 53;
    #10 ex_value = 11; ex_addr = 54;
    #10 ex_value = 230; ex_addr = 55;
    #10 ex_value = -40; ex_addr = 56;
    #10 ex_value = 190; ex_addr = 57;
    #10 ex_value = 47; ex_addr = 58;
    #10 ex_value = 251; ex_addr = 59;
    #10 ex_value = 249; ex_addr = 60;
    #10 ex_value = -90; ex_addr = 61;
    #10 ex_value = 239; ex_addr = 62;
    #10 ex_value = 38; ex_addr = 63;
    #10 ex_value = -254; ex_addr = 64;
    #10 ex_value = -155; ex_addr = 65;
    #10 ex_value = 63; ex_addr = 66;
    #10 ex_value = -55; ex_addr = 67;
    #10 ex_value = 161; ex_addr = 68;
    #10 ex_value = -237; ex_addr = 69;
    #10 ex_value = -50; ex_addr = 70;
    #10 ex_value = -120; ex_addr = 71;
    #10 ex_value = 138; ex_addr = 72;
    #10 ex_value = 66; ex_addr = 73;
    #10 ex_value = 66; ex_addr = 74;
    #10 ex_value = 103; ex_addr = 75;
    #10 ex_value = -236; ex_addr = 76;
    #10 ex_value = 238; ex_addr = 77;
    #10 ex_value = 38; ex_addr = 78;
    #10 ex_value = 244; ex_addr = 79;
    #10 ex_value = -88; ex_addr = 80;
    #10 ex_value = 120; ex_addr = 81;
    #10 ex_value = -61; ex_addr = 82;
    #10 ex_value = -160; ex_addr = 83;
    #10 ex_value = 149; ex_addr = 84;
    #10 ex_value = 104; ex_addr = 85;
    #10 ex_value = -246; ex_addr = 86;
    #10 ex_value = -82; ex_addr = 87;
    #10 ex_value = 181; ex_addr = 88;
    #10 ex_value = 216; ex_addr = 89;
    #10 ex_value = -108; ex_addr = 90;
    #10 ex_value = 207; ex_addr = 91;
    #10 ex_value = -135; ex_addr = 92;
    #10 ex_value = -171; ex_addr = 93;
    #10 ex_value = -161; ex_addr = 94;
    #10 ex_value = -114; ex_addr = 95;
    #10 ex_value = -239; ex_addr = 96;
    #10 ex_value = -222; ex_addr = 97;
    #10 ex_value = 93; ex_addr = 98;
    #10 ex_value = -62; ex_addr = 99;
    #10 ex_value = 177; ex_addr = 100;
    #10 ex_value = -186; ex_addr = 101;
    #10 ex_value = 217; ex_addr = 102;
    #10 ex_value = -120; ex_addr = 103;
    #10 ex_value = -224; ex_addr = 104;
    #10 ex_value = 213; ex_addr = 105;
    #10 ex_value = 220; ex_addr = 106;
    #10 ex_value = 117; ex_addr = 107;
    #10 ex_value = 67; ex_addr = 108;
    #10 ex_value = 179; ex_addr = 109;
    #10 ex_value = 200; ex_addr = 110;
    #10 ex_value = -166; ex_addr = 111;
    #10 ex_value = 57; ex_addr = 112;
    #10 ex_value = 232; ex_addr = 113;
    #10 ex_value = 69; ex_addr = 114;
    #10 ex_value = -36; ex_addr = 115;
    #10 ex_value = 223; ex_addr = 116;
    #10 ex_value = -211; ex_addr = 117;
    #10 ex_value = -209; ex_addr = 118;
    #10 ex_value = 164; ex_addr = 119;
    #10 ex_value = 104; ex_addr = 120;
    #10 ex_value = -150; ex_addr = 121;
    #10 ex_value = -225; ex_addr = 122;
    #10 ex_value = -85; ex_addr = 123;
    #10 ex_value = 239; ex_addr = 124;
    #10 ex_value = 67; ex_addr = 125;
    #10 ex_value = 247; ex_addr = 126;
    #10 ex_value = 154; ex_addr = 127;
    #10 ex_value = -124; ex_addr = 128;
    #10 ex_value = 129; ex_addr = 129;
    #10 ex_value = -207; ex_addr = 130;
    #10 ex_value = -28; ex_addr = 131;
    #10 ex_value = 135; ex_addr = 132;
    #10 ex_value = 73; ex_addr = 133;
    #10 ex_value = 181; ex_addr = 134;
    #10 ex_value = 87; ex_addr = 135;
    #10 ex_value = -169; ex_addr = 136;
    #10 ex_value = -174; ex_addr = 137;
    #10 ex_value = 147; ex_addr = 138;
    #10 ex_value = -54; ex_addr = 139;
    #10 ex_value = 254; ex_addr = 140;
    #10 ex_value = -177; ex_addr = 141;
    #10 ex_value = -142; ex_addr = 142;
    #10 ex_value = -213; ex_addr = 143;
    #10 ex_value = -7; ex_addr = 144;
    #10 ex_value = -120; ex_addr = 145;
    #10 ex_value = -250; ex_addr = 146;
    #10 ex_value = 10; ex_addr = 147;
    #10 ex_value = 63; ex_addr = 148;
    #10 ex_value = 2; ex_addr = 149;
    #10 ex_value = 234; ex_addr = 150;
    #10 ex_value = 9; ex_addr = 151;
    #10 ex_value = -242; ex_addr = 152;
    #10 ex_value = -173; ex_addr = 153;
    #10 ex_value = 161; ex_addr = 154;
    #10 ex_value = -29; ex_addr = 155;
    #10 ex_value = -23; ex_addr = 156;
    #10 ex_value = 193; ex_addr = 157;
    #10 ex_value = 232; ex_addr = 158;
    #10 ex_value = -180; ex_addr = 159;
    #10 ex_value = -38; ex_addr = 160;
    #10 ex_value = 36; ex_addr = 161;
    #10 ex_value = 108; ex_addr = 162;
    #10 ex_value = -179; ex_addr = 163;
    #10 ex_value = -168; ex_addr = 164;
    #10 ex_value = -47; ex_addr = 165;
    #10 ex_value = -36; ex_addr = 166;
    #10 ex_value = 18; ex_addr = 167;
    #10 ex_value = 24; ex_addr = 168;
    #10 ex_value = -36; ex_addr = 169;
    #10 ex_value = -67; ex_addr = 170;
    #10 ex_value = -208; ex_addr = 171;
    #10 ex_value = -176; ex_addr = 172;
    #10 ex_value = 99; ex_addr = 173;
    #10 ex_value = -43; ex_addr = 174;
    #10 ex_value = -157; ex_addr = 175;
    #10 ex_value = -6; ex_addr = 176;
    #10 ex_value = -145; ex_addr = 177;
    #10 ex_value = -138; ex_addr = 178;
    #10 ex_value = 214; ex_addr = 179;
    #10 ex_value = 15; ex_addr = 180;
    #10 ex_value = 224; ex_addr = 181;
    #10 ex_value = -25; ex_addr = 182;
    #10 ex_value = -149; ex_addr = 183;
    #10 ex_value = 171; ex_addr = 184;
    #10 ex_value = 68; ex_addr = 185;
    #10 ex_value = 135; ex_addr = 186;
    #10 ex_value = -99; ex_addr = 187;
    #10 ex_value = 120; ex_addr = 188;
    #10 ex_value = 226; ex_addr = 189;
    #10 ex_value = 99; ex_addr = 190;
    #10 ex_value = -216; ex_addr = 191;
    #10 ex_value = -169; ex_addr = 192;
    #10 ex_value = 118; ex_addr = 193;
    #10 ex_value = 34; ex_addr = 194;
    #10 ex_value = -186; ex_addr = 195;
    #10 ex_value = -46; ex_addr = 196;
    #10 ex_value = -25; ex_addr = 197;
    #10 ex_value = -130; ex_addr = 198;
    #10 ex_value = 82; ex_addr = 199;
    #10 ex_value = -129; ex_addr = 200;
    #10 ex_value = -219; ex_addr = 201;
    #10 ex_value = 229; ex_addr = 202;
    #10 ex_value = 8; ex_addr = 203;
    #10 ex_value = -224; ex_addr = 204;
    #10 ex_value = -134; ex_addr = 205;
    #10 ex_value = 198; ex_addr = 206;
    #10 ex_value = -210; ex_addr = 207;
    #10 ex_value = 173; ex_addr = 208;
    #10 ex_value = 15; ex_addr = 209;
    #10 ex_value = 27; ex_addr = 210;
    #10 ex_value = -80; ex_addr = 211;
    #10 ex_value = -193; ex_addr = 212;
    #10 ex_value = 190; ex_addr = 213;
    #10 ex_value = 56; ex_addr = 214;
    #10 ex_value = -109; ex_addr = 215;
    #10 ex_value = -126; ex_addr = 216;
    #10 ex_value = -159; ex_addr = 217;
    #10 ex_value = 141; ex_addr = 218;
    #10 ex_value = 234; ex_addr = 219;
    #10 WE = 1'b0;
    
    //first right answer
    //input right answer at ram2
    #10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b1;
    WE = 1'b1;
    #10 ex_value = 0; ex_addr = 10;
    #10 ex_value = 0; ex_addr = 11;
    #10 ex_value = 0; ex_addr = 12;
    #10 ex_value = 1536; ex_addr = 13;
    #10 ex_value = 0; ex_addr = 14;
    #10 ex_value = 0; ex_addr = 15;
    #10 ex_value = 0; ex_addr = 16;
    #10 ex_value = 0; ex_addr = 17;
    #10 ex_value = 0; ex_addr = 18;
    #10 ex_value = 0; ex_addr = 19;
    #10 WE = 1'b0;
    #10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b0;
    
	#10 ENABLE = 1'b1; WE = 1'b0;
	#20000;
    BCK_PROP_START = 1'b1; ENABLE = 1'b0;
    #20000;
    BCK_PROP_START = 1'b0;
    #10;
    
    //another right answer test bench - if need, make comment below section
    //---------------------------------------------------------------------
    //second right answer
    //input right answer at ram2
    /*#10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b1;
    for (i=0; i<BCK_CELL; i = i+1) begin
            ex_value = 0;
            WE = 1'b1;
            ex_addr = BCK_CELL + i;
            #10;
    end
    ex_addr = BCK_CELL + 1;
    ex_value = (1'b1 << 10) + (1'b1 << 9);
    #10 WE = 1'b0;
    #10 WEIGHT1 = 1'b0; WEIGHT2 = 1'b0; RIGHT_ANSWER = 1'b0;
    #10 ENABLE = 1'b1; WE = 1'b0;
	#5000;
    BCK_PROP_START = 1'b1; ENABLE = 1'b0;
    #3000;
    BCK_PROP_START = 1'b0;
    #10;*/
    //--------------------------------------------------------------------
    
    //BATCH_END = 1'b1;
    #5000;
    $stop;
end

endmodule