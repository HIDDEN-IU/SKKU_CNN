`timescale 1ns/1ns
module TOP_MODULE_CONV_tb(
);

reg CLK;
reg RESET_N;

reg [15:0] DATA, ADDR;
reg WE, CONV_WEIGHT1, CONV_WEIGHT2, CONV_WEIGHT3, IMG_INPUT,
    SRT_LAYER1, SRT_LAYER2, SRT_LAYER3;

wire DONE_LAYER1, DONE_LAYER2, DONE_LAYER3, WE_OUT;
wire [15:0] FLAT_OUT, ADDR_OUT;


integer signed i, j;

initial
begin
CLK = 0;
end

initial
begin
	forever
	begin
		#5 CLK = !CLK;
	end
end

TOP_MODULE_CONV top_module_conv(
.clk(CLK),
.reset_n(RESET_N),
.data(DATA),
.addr(ADDR),
.we(WE),
.conv_weight1(CONV_WEIGHT1),
.conv_weight2(CONV_WEIGHT2),
.conv_weight3(CONV_WEIGHT3),
.img_input(IMG_INPUT),
.srt_layer1(SRT_LAYER1),  //
.srt_layer2(SRT_LAYER2),  //
.srt_layer3(SRT_LAYER3),  //

.done_layer1(DONE_LAYER1),      //
.done_layer2(DONE_LAYER2),      //
.done_layer3(DONE_LAYER3),      //
.flat_out(FLAT_OUT),
.addr_out(ADDR_OUT),
.we_out(WE_OUT)
);

initial
begin
    {CONV_WEIGHT1, CONV_WEIGHT2, CONV_WEIGHT3, IMG_INPUT,
    SRT_LAYER1,SRT_LAYER2, SRT_LAYER3} <= 1'B0;
	RESET_N = 1'B0;
    #15 RESET_N = 1'B1;
    DATA = 1'B0; ADDR = 1'B0; WE = 1'b0;
    #10 CONV_WEIGHT1 = 1'B1;
    begin
    #10 DATA = -255; ADDR = 0; WE = 1'B1;
    #10 DATA = -255; ADDR = 1;
    #10 DATA = -255; ADDR = 2;
    #10 DATA = 0; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = 0; ADDR = 5;
    #10 DATA = 256; ADDR = 6;
    #10 DATA = 256; ADDR = 7;
    #10 DATA = 256; ADDR = 8;
    #10 DATA = 256; ADDR = 0;
    #10 DATA = 256; ADDR = 1;
    #10 DATA = 256; ADDR = 2;
    #10 DATA = 0; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = 0; ADDR = 5;
    #10 DATA = -255; ADDR = 6;
    #10 DATA = -255; ADDR = 7;
    #10 DATA = -255; ADDR = 8;
    #10 DATA = -255; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = 256; ADDR = 2;
    #10 DATA = -255; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = 256; ADDR = 5;
    #10 DATA = -255; ADDR = 6;
    #10 DATA = 0; ADDR = 7;
    #10 DATA = 256; ADDR = 8;
    #10 DATA = 256; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = -255; ADDR = 2;
    #10 DATA = 256; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = -255; ADDR = 5;
    #10 DATA = 256; ADDR = 6;
    #10 DATA = 0; ADDR = 7;
    #10 DATA = -255; ADDR = 8;
    #10 DATA = 256; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = -255; ADDR = 2;
    #10 DATA = 0; ADDR = 3;
    #10 DATA = 256; ADDR = 4;
    #10 DATA = 0; ADDR = 5;
    #10 DATA = -255; ADDR = 6;
    #10 DATA = 0; ADDR = 7;
    #10 DATA = 256; ADDR = 8;
    #10 DATA = -255; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = 256; ADDR = 2;
    #10 DATA = 0; ADDR = 3;
    #10 DATA = 256; ADDR = 4;
    #10 DATA = 0; ADDR = 5;
    #10 DATA = 256; ADDR = 6;
    #10 DATA = 0; ADDR = 7;
    #10 DATA = -255; ADDR = 8;
    end
    #20 WE = 1'b0;
    #10 CONV_WEIGHT1 = 1'B0;
    
    CONV_WEIGHT2 = 1'B1;
    begin
    #10 DATA = 23; ADDR = 0;WE = 1'B1;
    #10 DATA = -1; ADDR = 1;
    #10 DATA = 24; ADDR = 2;
    #10 DATA = 2; ADDR = 3;
    #10 DATA = 13; ADDR = 4;
    #10 DATA = 18; ADDR = 5;
    #10 DATA = -23; ADDR = 6;
    #10 DATA = 5; ADDR = 7;
    #10 DATA = 16; ADDR = 8;
    #10 DATA = 15; ADDR = 0;
    #10 DATA = 3; ADDR = 1;
    #10 DATA = 16; ADDR = 2;
    #10 DATA = -9; ADDR = 3;
    #10 DATA = -22; ADDR = 4;
    #10 DATA = 12; ADDR = 5;
    #10 DATA = -6; ADDR = 6;
    #10 DATA = 20; ADDR = 7;
    #10 DATA = 12; ADDR = 8;
    #10 DATA = -1; ADDR = 0;
    #10 DATA = -6; ADDR = 1;
    #10 DATA = -11; ADDR = 2;
    #10 DATA = -20; ADDR = 3;
    #10 DATA = -1; ADDR = 4;
    #10 DATA = 20; ADDR = 5;
    #10 DATA = 24; ADDR = 6;
    #10 DATA = 18; ADDR = 7;
    #10 DATA = 12; ADDR = 8;
    #10 DATA = 18; ADDR = 0;
    #10 DATA = -7; ADDR = 1;
    #10 DATA = -11; ADDR = 2;
    #10 DATA = -19; ADDR = 3;
    #10 DATA = 15; ADDR = 4;
    #10 DATA = -14; ADDR = 5;
    #10 DATA = 22; ADDR = 6;
    #10 DATA = 3; ADDR = 7;
    #10 DATA = 6; ADDR = 8;
    #10 DATA = -13; ADDR = 0;
    #10 DATA = 15; ADDR = 1;
    #10 DATA = -13; ADDR = 2;
    #10 DATA = -5; ADDR = 3;
    #10 DATA = 18; ADDR = 4;
    #10 DATA = -16; ADDR = 5;
    #10 DATA = -13; ADDR = 6;
    #10 DATA = -1; ADDR = 7;
    #10 DATA = 14; ADDR = 8;
    #10 DATA = 1; ADDR = 0;
    #10 DATA = 5; ADDR = 1;
    #10 DATA = 0; ADDR = 2;
    #10 DATA = -25; ADDR = 3;
    #10 DATA = -9; ADDR = 4;
    #10 DATA = 6; ADDR = 5;
    #10 DATA = 0; ADDR = 6;
    #10 DATA = -21; ADDR = 7;
    #10 DATA = 0; ADDR = 8;
    #10 DATA = -21; ADDR = 0;
    #10 DATA = -9; ADDR = 1;
    #10 DATA = 16; ADDR = 2;
    #10 DATA = 16; ADDR = 3;
    #10 DATA = -5; ADDR = 4;
    #10 DATA = -10; ADDR = 5;
    #10 DATA = 23; ADDR = 6;
    #10 DATA = 24; ADDR = 7;
    #10 DATA = 13; ADDR = 8;
    #10 DATA = 5; ADDR = 0;
    #10 DATA = 19; ADDR = 1;
    #10 DATA = -22; ADDR = 2;
    #10 DATA = -10; ADDR = 3;
    #10 DATA = -8; ADDR = 4;
    #10 DATA = -15; ADDR = 5;
    #10 DATA = 12; ADDR = 6;
    #10 DATA = 23; ADDR = 7;
    #10 DATA = 9; ADDR = 8;
    #10 DATA = 13; ADDR = 0;
    #10 DATA = 19; ADDR = 1;
    #10 DATA = 1; ADDR = 2;
    #10 DATA = -3; ADDR = 3;
    #10 DATA = 13; ADDR = 4;
    #10 DATA = 25; ADDR = 5;
    #10 DATA = -18; ADDR = 6;
    #10 DATA = -19; ADDR = 7;
    #10 DATA = 0; ADDR = 8;
    #10 DATA = 15; ADDR = 0;
    #10 DATA = 23; ADDR = 1;
    #10 DATA = 22; ADDR = 2;
    #10 DATA = 9; ADDR = 3;
    #10 DATA = -2; ADDR = 4;
    #10 DATA = 20; ADDR = 5;
    #10 DATA = 4; ADDR = 6;
    #10 DATA = -12; ADDR = 7;
    #10 DATA = -22; ADDR = 8;
    #10 DATA = 18; ADDR = 0;
    #10 DATA = 5; ADDR = 1;
    #10 DATA = 12; ADDR = 2;
    #10 DATA = 12; ADDR = 3;
    #10 DATA = 15; ADDR = 4;
    #10 DATA = 8; ADDR = 5;
    #10 DATA = -13; ADDR = 6;
    #10 DATA = -17; ADDR = 7;
    #10 DATA = 1; ADDR = 8;
    #10 DATA = -6; ADDR = 0;
    #10 DATA = -21; ADDR = 1;
    #10 DATA = 24; ADDR = 2;
    #10 DATA = -13; ADDR = 3;
    #10 DATA = -24; ADDR = 4;
    #10 DATA = 15; ADDR = 5;
    #10 DATA = -22; ADDR = 6;
    #10 DATA = 14; ADDR = 7;
    #10 DATA = 20; ADDR = 8;
    #10 DATA = -20; ADDR = 0;
    #10 DATA = 18; ADDR = 1;
    #10 DATA = -21; ADDR = 2;
    #10 DATA = 15; ADDR = 3;
    #10 DATA = 24; ADDR = 4;
    #10 DATA = 4; ADDR = 5;
    #10 DATA = -5; ADDR = 6;
    #10 DATA = -8; ADDR = 7;
    #10 DATA = 9; ADDR = 8;
    #10 DATA = 25; ADDR = 0;
    #10 DATA = -7; ADDR = 1;
    #10 DATA = -13; ADDR = 2;
    #10 DATA = 19; ADDR = 3;
    #10 DATA = -7; ADDR = 4;
    #10 DATA = 10; ADDR = 5;
    #10 DATA = -7; ADDR = 6;
    #10 DATA = 7; ADDR = 7;
    #10 DATA = 1; ADDR = 8;
    #10 DATA = 12; ADDR = 0;
    #10 DATA = -19; ADDR = 1;
    #10 DATA = -2; ADDR = 2;
    #10 DATA = 3; ADDR = 3;
    #10 DATA = -4; ADDR = 4;
    #10 DATA = -25; ADDR = 5;
    #10 DATA = -12; ADDR = 6;
    #10 DATA = 13; ADDR = 7;
    #10 DATA = 5; ADDR = 8;
    #10 DATA = 17; ADDR = 0;
    #10 DATA = 7; ADDR = 1;
    #10 DATA = 11; ADDR = 2;
    #10 DATA = 4; ADDR = 3;
    #10 DATA = -11; ADDR = 4;
    #10 DATA = -13; ADDR = 5;
    #10 DATA = -23; ADDR = 6;
    #10 DATA = -8; ADDR = 7;
    #10 DATA = -13; ADDR = 8;
    end
    #20 WE = 1'b0;
    #10 CONV_WEIGHT2 = 1'B0;
    
    CONV_WEIGHT3 = 1'B1;
    begin
    #10 DATA = -22; ADDR = 0;WE = 1'B1;
    #10 DATA = -21; ADDR = 1;
    #10 DATA = 5; ADDR = 2;
    #10 DATA = 13; ADDR = 3;
    #10 DATA = 8; ADDR = 4;
    #10 DATA = -17; ADDR = 5;
    #10 DATA = 11; ADDR = 6;
    #10 DATA = 13; ADDR = 7;
    #10 DATA = -19; ADDR = 8;
    #10 DATA = 8; ADDR = 0;
    #10 DATA = 10; ADDR = 1;
    #10 DATA = -23; ADDR = 2;
    #10 DATA = -13; ADDR = 3;
    #10 DATA = -5; ADDR = 4;
    #10 DATA = -12; ADDR = 5;
    #10 DATA = 22; ADDR = 6;
    #10 DATA = -9; ADDR = 7;
    #10 DATA = -4; ADDR = 8;
    #10 DATA = 10; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = -1; ADDR = 2;
    #10 DATA = -8; ADDR = 3;
    #10 DATA = 14; ADDR = 4;
    #10 DATA = -5; ADDR = 5;
    #10 DATA = -4; ADDR = 6;
    #10 DATA = -12; ADDR = 7;
    #10 DATA = 16; ADDR = 8;
    #10 DATA = -23; ADDR = 0;
    #10 DATA = 3; ADDR = 1;
    #10 DATA = -2; ADDR = 2;
    #10 DATA = -17; ADDR = 3;
    #10 DATA = -12; ADDR = 4;
    #10 DATA = 23; ADDR = 5;
    #10 DATA = 3; ADDR = 6;
    #10 DATA = -15; ADDR = 7;
    #10 DATA = 24; ADDR = 8;
    #10 DATA = -24; ADDR = 0;
    #10 DATA = -8; ADDR = 1;
    #10 DATA = 19; ADDR = 2;
    #10 DATA = 13; ADDR = 3;
    #10 DATA = 22; ADDR = 4;
    #10 DATA = -18; ADDR = 5;
    #10 DATA = 15; ADDR = 6;
    #10 DATA = 25; ADDR = 7;
    #10 DATA = 12; ADDR = 8;
    #10 DATA = 20; ADDR = 0;
    #10 DATA = -18; ADDR = 1;
    #10 DATA = -11; ADDR = 2;
    #10 DATA = 5; ADDR = 3;
    #10 DATA = -16; ADDR = 4;
    #10 DATA = 8; ADDR = 5;
    #10 DATA = -3; ADDR = 6;
    #10 DATA = -11; ADDR = 7;
    #10 DATA = -20; ADDR = 8;
    #10 DATA = 3; ADDR = 0;
    #10 DATA = 13; ADDR = 1;
    #10 DATA = 24; ADDR = 2;
    #10 DATA = 13; ADDR = 3;
    #10 DATA = 2; ADDR = 4;
    #10 DATA = 20; ADDR = 5;
    #10 DATA = 12; ADDR = 6;
    #10 DATA = 7; ADDR = 7;
    #10 DATA = 24; ADDR = 8;
    #10 DATA = -23; ADDR = 0;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = -10; ADDR = 2;
    #10 DATA = 20; ADDR = 3;
    #10 DATA = 19; ADDR = 4;
    #10 DATA = 12; ADDR = 5;
    #10 DATA = -19; ADDR = 6;
    #10 DATA = -14; ADDR = 7;
    #10 DATA = -13; ADDR = 8;
    #10 DATA = -23; ADDR = 0;
    #10 DATA = 15; ADDR = 1;
    #10 DATA = -21; ADDR = 2;
    #10 DATA = -7; ADDR = 3;
    #10 DATA = 24; ADDR = 4;
    #10 DATA = -2; ADDR = 5;
    #10 DATA = 7; ADDR = 6;
    #10 DATA = -4; ADDR = 7;
    #10 DATA = -19; ADDR = 8;
    #10 DATA = 22; ADDR = 0;
    #10 DATA = -22; ADDR = 1;
    #10 DATA = -14; ADDR = 2;
    #10 DATA = 15; ADDR = 3;
    #10 DATA = 17; ADDR = 4;
    #10 DATA = -24; ADDR = 5;
    #10 DATA = 0; ADDR = 6;
    #10 DATA = -12; ADDR = 7;
    #10 DATA = 16; ADDR = 8;
    #10 DATA = -25; ADDR = 0;
    #10 DATA = 6; ADDR = 1;
    #10 DATA = -5; ADDR = 2;
    #10 DATA = -22; ADDR = 3;
    #10 DATA = -8; ADDR = 4;
    #10 DATA = 8; ADDR = 5;
    #10 DATA = 16; ADDR = 6;
    #10 DATA = 8; ADDR = 7;
    #10 DATA = 22; ADDR = 8;
    #10 DATA = 7; ADDR = 0;
    #10 DATA = 1; ADDR = 1;
    #10 DATA = -16; ADDR = 2;
    #10 DATA = -6; ADDR = 3;
    #10 DATA = -1; ADDR = 4;
    #10 DATA = 17; ADDR = 5;
    #10 DATA = -19; ADDR = 6;
    #10 DATA = 1; ADDR = 7;
    #10 DATA = 14; ADDR = 8;
    #10 DATA = -25; ADDR = 0;
    #10 DATA = -17; ADDR = 1;
    #10 DATA = 6; ADDR = 2;
    #10 DATA = 4; ADDR = 3;
    #10 DATA = -25; ADDR = 4;
    #10 DATA = -3; ADDR = 5;
    #10 DATA = 25; ADDR = 6;
    #10 DATA = 21; ADDR = 7;
    #10 DATA = -10; ADDR = 8;
    #10 DATA = 21; ADDR = 0;
    #10 DATA = 18; ADDR = 1;
    #10 DATA = -13; ADDR = 2;
    #10 DATA = -2; ADDR = 3;
    #10 DATA = 19; ADDR = 4;
    #10 DATA = 10; ADDR = 5;
    #10 DATA = -6; ADDR = 6;
    #10 DATA = -20; ADDR = 7;
    #10 DATA = -1; ADDR = 8;
    #10 DATA = -8; ADDR = 0;
    #10 DATA = 3; ADDR = 1;
    #10 DATA = 14; ADDR = 2;
    #10 DATA = 11; ADDR = 3;
    #10 DATA = -4; ADDR = 4;
    #10 DATA = 12; ADDR = 5;
    #10 DATA = 11; ADDR = 6;
    #10 DATA = -11; ADDR = 7;
    #10 DATA = -2; ADDR = 8;
    #10 DATA = 6; ADDR = 0;
    #10 DATA = -11; ADDR = 1;
    #10 DATA = -20; ADDR = 2;
    #10 DATA = 7; ADDR = 3;
    #10 DATA = 4; ADDR = 4;
    #10 DATA = 4; ADDR = 5;
    #10 DATA = 8; ADDR = 6;
    #10 DATA = -21; ADDR = 7;
    #10 DATA = -6; ADDR = 8;
    #10 DATA = -15; ADDR = 0;
    #10 DATA = -9; ADDR = 1;
    #10 DATA = -2; ADDR = 2;
    #10 DATA = 15; ADDR = 3;
    #10 DATA = -8; ADDR = 4;
    #10 DATA = -1; ADDR = 5;
    #10 DATA = 16; ADDR = 6;
    #10 DATA = 20; ADDR = 7;
    #10 DATA = 3; ADDR = 8;
    #10 DATA = -21; ADDR = 0;
    #10 DATA = 4; ADDR = 1;
    #10 DATA = 3; ADDR = 2;
    #10 DATA = -14; ADDR = 3;
    #10 DATA = 4; ADDR = 4;
    #10 DATA = -10; ADDR = 5;
    #10 DATA = -16; ADDR = 6;
    #10 DATA = -8; ADDR = 7;
    #10 DATA = -24; ADDR = 8;
    #10 DATA = 20; ADDR = 0;
    #10 DATA = -23; ADDR = 1;
    #10 DATA = 19; ADDR = 2;
    #10 DATA = -22; ADDR = 3;
    #10 DATA = -8; ADDR = 4;
    #10 DATA = 14; ADDR = 5;
    #10 DATA = -4; ADDR = 6;
    #10 DATA = -4; ADDR = 7;
    #10 DATA = 25; ADDR = 8;
    #10 DATA = 14; ADDR = 0;
    #10 DATA = 18; ADDR = 1;
    #10 DATA = -19; ADDR = 2;
    #10 DATA = -25; ADDR = 3;
    #10 DATA = -4; ADDR = 4;
    #10 DATA = -20; ADDR = 5;
    #10 DATA = -15; ADDR = 6;
    #10 DATA = 22; ADDR = 7;
    #10 DATA = 17; ADDR = 8;
    #10 DATA = 24; ADDR = 0;
    #10 DATA = 17; ADDR = 1;
    #10 DATA = 5; ADDR = 2;
    #10 DATA = 23; ADDR = 3;
    #10 DATA = -17; ADDR = 4;
    #10 DATA = -5; ADDR = 5;
    #10 DATA = 6; ADDR = 6;
    #10 DATA = 18; ADDR = 7;
    #10 DATA = 25; ADDR = 8;
    #10 DATA = -13; ADDR = 0;
    #10 DATA = -4; ADDR = 1;
    #10 DATA = 15; ADDR = 2;
    #10 DATA = 20; ADDR = 3;
    #10 DATA = 8; ADDR = 4;
    #10 DATA = -10; ADDR = 5;
    #10 DATA = -19; ADDR = 6;
    #10 DATA = -7; ADDR = 7;
    #10 DATA = 17; ADDR = 8;
    #10 DATA = -12; ADDR = 0;
    #10 DATA = 9; ADDR = 1;
    #10 DATA = 21; ADDR = 2;
    #10 DATA = 22; ADDR = 3;
    #10 DATA = 17; ADDR = 4;
    #10 DATA = 13; ADDR = 5;
    #10 DATA = -14; ADDR = 6;
    #10 DATA = -3; ADDR = 7;
    #10 DATA = -19; ADDR = 8;
    #10 DATA = -1; ADDR = 0;
    #10 DATA = 22; ADDR = 1;
    #10 DATA = 23; ADDR = 2;
    #10 DATA = -22; ADDR = 3;
    #10 DATA = -25; ADDR = 4;
    #10 DATA = -25; ADDR = 5;
    #10 DATA = 6; ADDR = 6;
    #10 DATA = -19; ADDR = 7;
    #10 DATA = 15; ADDR = 8;
    #10 DATA = -10; ADDR = 0;
    #10 DATA = 18; ADDR = 1;
    #10 DATA = 1; ADDR = 2;
    #10 DATA = -19; ADDR = 3;
    #10 DATA = -12; ADDR = 4;
    #10 DATA = -22; ADDR = 5;
    #10 DATA = 2; ADDR = 6;
    #10 DATA = -9; ADDR = 7;
    #10 DATA = 18; ADDR = 8;
    #10 DATA = -24; ADDR = 0;
    #10 DATA = -7; ADDR = 1;
    #10 DATA = 17; ADDR = 2;
    #10 DATA = 14; ADDR = 3;
    #10 DATA = 11; ADDR = 4;
    #10 DATA = 7; ADDR = 5;
    #10 DATA = -6; ADDR = 6;
    #10 DATA = -4; ADDR = 7;
    #10 DATA = -25; ADDR = 8;
    #10 DATA = 8; ADDR = 0;
    #10 DATA = -2; ADDR = 1;
    #10 DATA = 8; ADDR = 2;
    #10 DATA = 4; ADDR = 3;
    #10 DATA = -19; ADDR = 4;
    #10 DATA = 6; ADDR = 5;
    #10 DATA = -14; ADDR = 6;
    #10 DATA = 3; ADDR = 7;
    #10 DATA = -7; ADDR = 8;
    #10 DATA = 0; ADDR = 0;
    #10 DATA = -4; ADDR = 1;
    #10 DATA = 24; ADDR = 2;
    #10 DATA = -2; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = -12; ADDR = 5;
    #10 DATA = 22; ADDR = 6;
    #10 DATA = 2; ADDR = 7;
    #10 DATA = -20; ADDR = 8;
    #10 DATA = 20; ADDR = 0;
    #10 DATA = -10; ADDR = 1;
    #10 DATA = -15; ADDR = 2;
    #10 DATA = -19; ADDR = 3;
    #10 DATA = -18; ADDR = 4;
    #10 DATA = 6; ADDR = 5;
    #10 DATA = -6; ADDR = 6;
    #10 DATA = -7; ADDR = 7;
    #10 DATA = 11; ADDR = 8;
    #10 DATA = 19; ADDR = 0;
    #10 DATA = -8; ADDR = 1;
    #10 DATA = -7; ADDR = 2;
    #10 DATA = -17; ADDR = 3;
    #10 DATA = 17; ADDR = 4;
    #10 DATA = 23; ADDR = 5;
    #10 DATA = 25; ADDR = 6;
    #10 DATA = 23; ADDR = 7;
    #10 DATA = -6; ADDR = 8;
    #10 DATA = -14; ADDR = 0;
    #10 DATA = -22; ADDR = 1;
    #10 DATA = 10; ADDR = 2;
    #10 DATA = 8; ADDR = 3;
    #10 DATA = -21; ADDR = 4;
    #10 DATA = 12; ADDR = 5;
    #10 DATA = -10; ADDR = 6;
    #10 DATA = 11; ADDR = 7;
    #10 DATA = 7; ADDR = 8;
    #10 DATA = -5; ADDR = 0;
    #10 DATA = 1; ADDR = 1;
    #10 DATA = 7; ADDR = 2;
    #10 DATA = 21; ADDR = 3;
    #10 DATA = -23; ADDR = 4;
    #10 DATA = 5; ADDR = 5;
    #10 DATA = -13; ADDR = 6;
    #10 DATA = -13; ADDR = 7;
    #10 DATA = -5; ADDR = 8;
    end
    #20 WE = 1'B0;
    #10 CONV_WEIGHT3 = 1'B0; 
    
    IMG_INPUT = 1'B1;
    begin
    #10 DATA = 0; ADDR = 0; WE = 1'b1;
    #10 DATA = 0; ADDR = 1;
    #10 DATA = 0; ADDR = 2;
    #10 DATA = 0; ADDR = 3;
    #10 DATA = 0; ADDR = 4;
    #10 DATA = 0; ADDR = 5;
    #10 DATA = 0; ADDR = 6;
    #10 DATA = 0; ADDR = 7;
    #10 DATA = 0; ADDR = 8;
    #10 DATA = 0; ADDR = 9;
    #10 DATA = 0; ADDR = 10;
    #10 DATA = 0; ADDR = 11;
    #10 DATA = 0; ADDR = 12;
    #10 DATA = 0; ADDR = 13;
    #10 DATA = 0; ADDR = 14;
    #10 DATA = 0; ADDR = 15;
    #10 DATA = 0; ADDR = 16;
    #10 DATA = 0; ADDR = 17;
    #10 DATA = 0; ADDR = 18;
    #10 DATA = 0; ADDR = 19;
    #10 DATA = 0; ADDR = 20;
    #10 DATA = 0; ADDR = 21;
    #10 DATA = 0; ADDR = 22;
    #10 DATA = 0; ADDR = 23;
    #10 DATA = 0; ADDR = 24;
    #10 DATA = 0; ADDR = 25;
    #10 DATA = 0; ADDR = 26;
    #10 DATA = 0; ADDR = 27;
    #10 DATA = 0; ADDR = 28;
    #10 DATA = 0; ADDR = 29;
    #10 DATA = 0; ADDR = 30;
    #10 DATA = 0; ADDR = 31;
    #10 DATA = 0; ADDR = 32;
    #10 DATA = 0; ADDR = 33;
    #10 DATA = 0; ADDR = 34;
    #10 DATA = 0; ADDR = 35;
    #10 DATA = 0; ADDR = 36;
    #10 DATA = 0; ADDR = 37;
    #10 DATA = 0; ADDR = 38;
    #10 DATA = 0; ADDR = 39;
    #10 DATA = 0; ADDR = 40;
    #10 DATA = 0; ADDR = 41;
    #10 DATA = 120; ADDR = 42;
    #10 DATA = 200; ADDR = 43;
    #10 DATA = 200; ADDR = 44;
    #10 DATA = 120; ADDR = 45;
    #10 DATA = 50; ADDR = 46;
    #10 DATA = 0; ADDR = 47;
    #10 DATA = 0; ADDR = 48;
    #10 DATA = 0; ADDR = 49;
    #10 DATA = 0; ADDR = 50;
    #10 DATA = 0; ADDR = 51;
    #10 DATA = 0; ADDR = 52;
    #10 DATA = 0; ADDR = 53;
    #10 DATA = 0; ADDR = 54;
    #10 DATA = 0; ADDR = 55;
    #10 DATA = 0; ADDR = 56;
    #10 DATA = 0; ADDR = 57;
    #10 DATA = 0; ADDR = 58;
    #10 DATA = 200; ADDR = 59;
    #10 DATA = 256; ADDR = 60;
    #10 DATA = 256; ADDR = 61;
    #10 DATA = 256; ADDR = 62;
    #10 DATA = 256; ADDR = 63;
    #10 DATA = 256; ADDR = 64;
    #10 DATA = 200; ADDR = 65;
    #10 DATA = 50; ADDR = 66;
    #10 DATA = 0; ADDR = 67;
    #10 DATA = 0; ADDR = 68;
    #10 DATA = 0; ADDR = 69;
    #10 DATA = 0; ADDR = 70;
    #10 DATA = 0; ADDR = 71;
    #10 DATA = 0; ADDR = 72;
    #10 DATA = 0; ADDR = 73;
    #10 DATA = 0; ADDR = 74;
    #10 DATA = 50; ADDR = 75;
    #10 DATA = 200; ADDR = 76;
    #10 DATA = 256; ADDR = 77;
    #10 DATA = 256; ADDR = 78;
    #10 DATA = 200; ADDR = 79;
    #10 DATA = 0; ADDR = 80;
    #10 DATA = 200; ADDR = 81;
    #10 DATA = 256; ADDR = 82;
    #10 DATA = 256; ADDR = 83;
    #10 DATA = 256; ADDR = 84;
    #10 DATA = 0; ADDR = 85;
    #10 DATA = 0; ADDR = 86;
    #10 DATA = 0; ADDR = 87;
    #10 DATA = 0; ADDR = 88;
    #10 DATA = 0; ADDR = 89;
    #10 DATA = 0; ADDR = 90;
    #10 DATA = 0; ADDR = 91;
    #10 DATA = 0; ADDR = 92;
    #10 DATA = 200; ADDR = 93;
    #10 DATA = 256; ADDR = 94;
    #10 DATA = 120; ADDR = 95;
    #10 DATA = 0; ADDR = 96;
    #10 DATA = 0; ADDR = 97;
    #10 DATA = 0; ADDR = 98;
    #10 DATA = 0; ADDR = 99;
    #10 DATA = 50; ADDR = 100;
    #10 DATA = 200; ADDR = 101;
    #10 DATA = 256; ADDR = 102;
    #10 DATA = 0; ADDR = 103;
    #10 DATA = 0; ADDR = 104;
    #10 DATA = 0; ADDR = 105;
    #10 DATA = 0; ADDR = 106;
    #10 DATA = 0; ADDR = 107;
    #10 DATA = 0; ADDR = 108;
    #10 DATA = 0; ADDR = 109;
    #10 DATA = 120; ADDR = 110;
    #10 DATA = 256; ADDR = 111;
    #10 DATA = 120; ADDR = 112;
    #10 DATA = 0; ADDR = 113;
    #10 DATA = 0; ADDR = 114;
    #10 DATA = 0; ADDR = 115;
    #10 DATA = 0; ADDR = 116;
    #10 DATA = 0; ADDR = 117;
    #10 DATA = 120; ADDR = 118;
    #10 DATA = 256; ADDR = 119;
    #10 DATA = 200; ADDR = 120;
    #10 DATA = 0; ADDR = 121;
    #10 DATA = 0; ADDR = 122;
    #10 DATA = 0; ADDR = 123;
    #10 DATA = 0; ADDR = 124;
    #10 DATA = 0; ADDR = 125;
    #10 DATA = 0; ADDR = 126;
    #10 DATA = 0; ADDR = 127;
    #10 DATA = 50; ADDR = 128;
    #10 DATA = 120; ADDR = 129;
    #10 DATA = 0; ADDR = 130;
    #10 DATA = 0; ADDR = 131;
    #10 DATA = 0; ADDR = 132;
    #10 DATA = 0; ADDR = 133;
    #10 DATA = 120; ADDR = 134;
    #10 DATA = 200; ADDR = 135;
    #10 DATA = 256; ADDR = 136;
    #10 DATA = 256; ADDR = 137;
    #10 DATA = 200; ADDR = 138;
    #10 DATA = 0; ADDR = 139;
    #10 DATA = 0; ADDR = 140;
    #10 DATA = 0; ADDR = 141;
    #10 DATA = 0; ADDR = 142;
    #10 DATA = 0; ADDR = 143;
    #10 DATA = 0; ADDR = 144;
    #10 DATA = 0; ADDR = 145;
    #10 DATA = 0; ADDR = 146;
    #10 DATA = 0; ADDR = 147;
    #10 DATA = 0; ADDR = 148;
    #10 DATA = 0; ADDR = 149;
    #10 DATA = 0; ADDR = 150;
    #10 DATA = 200; ADDR = 151;
    #10 DATA = 256; ADDR = 152;
    #10 DATA = 256; ADDR = 153;
    #10 DATA = 256; ADDR = 154;
    #10 DATA = 256; ADDR = 155;
    #10 DATA = 256; ADDR = 156;
    #10 DATA = 50; ADDR = 157;
    #10 DATA = 0; ADDR = 158;
    #10 DATA = 0; ADDR = 159;
    #10 DATA = 0; ADDR = 160;
    #10 DATA = 0; ADDR = 161;
    #10 DATA = 0; ADDR = 162;
    #10 DATA = 0; ADDR = 163;
    #10 DATA = 0; ADDR = 164;
    #10 DATA = 0; ADDR = 165;
    #10 DATA = 0; ADDR = 166;
    #10 DATA = 0; ADDR = 167;
    #10 DATA = 200; ADDR = 168;
    #10 DATA = 256; ADDR = 169;
    #10 DATA = 200; ADDR = 170;
    #10 DATA = 120; ADDR = 171;
    #10 DATA = 50; ADDR = 172;
    #10 DATA = 200; ADDR = 173;
    #10 DATA = 256; ADDR = 174;
    #10 DATA = 200; ADDR = 175;
    #10 DATA = 0; ADDR = 176;
    #10 DATA = 0; ADDR = 177;
    #10 DATA = 0; ADDR = 178;
    #10 DATA = 0; ADDR = 179;
    #10 DATA = 0; ADDR = 180;
    #10 DATA = 0; ADDR = 181;
    #10 DATA = 0; ADDR = 182;
    #10 DATA = 0; ADDR = 183;
    #10 DATA = 0; ADDR = 184;
    #10 DATA = 120; ADDR = 185;
    #10 DATA = 256; ADDR = 186;
    #10 DATA = 200; ADDR = 187;
    #10 DATA = 0; ADDR = 188;
    #10 DATA = 0; ADDR = 189;
    #10 DATA = 0; ADDR = 190;
    #10 DATA = 120; ADDR = 191;
    #10 DATA = 256; ADDR = 192;
    #10 DATA = 256; ADDR = 193;
    #10 DATA = 0; ADDR = 194;
    #10 DATA = 0; ADDR = 195;
    #10 DATA = 0; ADDR = 196;
    #10 DATA = 0; ADDR = 197;
    #10 DATA = 0; ADDR = 198;
    #10 DATA = 0; ADDR = 199;
    #10 DATA = 0; ADDR = 200;
    #10 DATA = 0; ADDR = 201;
    #10 DATA = 0; ADDR = 202;
    #10 DATA = 50; ADDR = 203;
    #10 DATA = 120; ADDR = 204;
    #10 DATA = 0; ADDR = 205;
    #10 DATA = 0; ADDR = 206;
    #10 DATA = 0; ADDR = 207;
    #10 DATA = 0; ADDR = 208;
    #10 DATA = 200; ADDR = 209;
    #10 DATA = 256; ADDR = 210;
    #10 DATA = 256; ADDR = 211;
    #10 DATA = 0; ADDR = 212;
    #10 DATA = 0; ADDR = 213;
    #10 DATA = 0; ADDR = 214;
    #10 DATA = 0; ADDR = 215;
    #10 DATA = 0; ADDR = 216;
    #10 DATA = 0; ADDR = 217;
    #10 DATA = 0; ADDR = 218;
    #10 DATA = 0; ADDR = 219;
    #10 DATA = 0; ADDR = 220;
    #10 DATA = 0; ADDR = 221;
    #10 DATA = 0; ADDR = 222;
    #10 DATA = 0; ADDR = 223;
    #10 DATA = 0; ADDR = 224;
    #10 DATA = 0; ADDR = 225;
    #10 DATA = 200; ADDR = 226;
    #10 DATA = 256; ADDR = 227;
    #10 DATA = 256; ADDR = 228;
    #10 DATA = 120; ADDR = 229;
    #10 DATA = 0; ADDR = 230;
    #10 DATA = 0; ADDR = 231;
    #10 DATA = 0; ADDR = 232;
    #10 DATA = 0; ADDR = 233;
    #10 DATA = 0; ADDR = 234;
    #10 DATA = 0; ADDR = 235;
    #10 DATA = 0; ADDR = 236;
    #10 DATA = 0; ADDR = 237;
    #10 DATA = 0; ADDR = 238;
    #10 DATA = 0; ADDR = 239;
    #10 DATA = 0; ADDR = 240;
    #10 DATA = 0; ADDR = 241;
    #10 DATA = 200; ADDR = 242;
    #10 DATA = 256; ADDR = 243;
    #10 DATA = 256; ADDR = 244;
    #10 DATA = 200; ADDR = 245;
    #10 DATA = 120; ADDR = 246;
    #10 DATA = 0; ADDR = 247;
    #10 DATA = 0; ADDR = 248;
    #10 DATA = 0; ADDR = 249;
    #10 DATA = 0; ADDR = 250;
    #10 DATA = 0; ADDR = 251;
    #10 DATA = 0; ADDR = 252;
    #10 DATA = 0; ADDR = 253;
    #10 DATA = 0; ADDR = 254;
    #10 DATA = 0; ADDR = 255;
    #10 DATA = 0; ADDR = 256;
    #10 DATA = 0; ADDR = 257;
    #10 DATA = 0; ADDR = 258;
    #10 DATA = 200; ADDR = 259;
    #10 DATA = 256; ADDR = 260;
    #10 DATA = 256; ADDR = 261;
    #10 DATA = 200; ADDR = 262;
    #10 DATA = 50; ADDR = 263;
    #10 DATA = 0; ADDR = 264;
    #10 DATA = 0; ADDR = 265;
    #10 DATA = 0; ADDR = 266;
    #10 DATA = 0; ADDR = 267;
    #10 DATA = 0; ADDR = 268;
    #10 DATA = 0; ADDR = 269;
    #10 DATA = 0; ADDR = 270;
    #10 DATA = 0; ADDR = 271;
    #10 DATA = 0; ADDR = 272;
    #10 DATA = 0; ADDR = 273;
    #10 DATA = 0; ADDR = 274;
    #10 DATA = 0; ADDR = 275;
    #10 DATA = 120; ADDR = 276;
    #10 DATA = 256; ADDR = 277;
    #10 DATA = 200; ADDR = 278;
    #10 DATA = 120; ADDR = 279;
    #10 DATA = 0; ADDR = 280;
    #10 DATA = 0; ADDR = 281;
    #10 DATA = 0; ADDR = 282;
    #10 DATA = 0; ADDR = 283;
    #10 DATA = 0; ADDR = 284;
    #10 DATA = 0; ADDR = 285;
    #10 DATA = 0; ADDR = 286;
    #10 DATA = 0; ADDR = 287;
    #10 DATA = 0; ADDR = 288;
    #10 DATA = 0; ADDR = 289;
    #10 DATA = 0; ADDR = 290;
    #10 DATA = 0; ADDR = 291;
    #10 DATA = 0; ADDR = 292;
    #10 DATA = 0; ADDR = 293;
    #10 DATA = 50; ADDR = 294;
    #10 DATA = 50; ADDR = 295;
    #10 DATA = 50; ADDR = 296;
    #10 DATA = 0; ADDR = 297;
    #10 DATA = 0; ADDR = 298;
    #10 DATA = 0; ADDR = 299;
    #10 DATA = 0; ADDR = 300;
    #10 DATA = 0; ADDR = 301;
    #10 DATA = 0; ADDR = 302;
    #10 DATA = 0; ADDR = 303;
    #10 DATA = 0; ADDR = 304;
    #10 DATA = 0; ADDR = 305;
    #10 DATA = 0; ADDR = 306;
    #10 DATA = 0; ADDR = 307;
    #10 DATA = 0; ADDR = 308;
    #10 DATA = 0; ADDR = 309;
    #10 DATA = 0; ADDR = 310;
    #10 DATA = 0; ADDR = 311;
    #10 DATA = 0; ADDR = 312;
    #10 DATA = 0; ADDR = 313;
    #10 DATA = 0; ADDR = 314;
    #10 DATA = 0; ADDR = 315;
    #10 DATA = 0; ADDR = 316;
    #10 DATA = 0; ADDR = 317;
    #10 DATA = 0; ADDR = 318;
    #10 DATA = 0; ADDR = 319;
    #10 DATA = 0; ADDR = 320;
    #10 DATA = 0; ADDR = 321;
    #10 DATA = 0; ADDR = 322;
    #10 DATA = 0; ADDR = 323;
    end
    #20 WE = 1'b0; 
    #10 IMG_INPUT = 1'B0;
    SRT_LAYER1 = 1'B1;
    wait(DONE_LAYER1); SRT_LAYER1 = 1'B0; SRT_LAYER2 = 1'B1; $stop; 
    wait(DONE_LAYER2); SRT_LAYER2 = 1'B0; SRT_LAYER3 = 1'B1; $stop; 
    wait(DONE_LAYER3); SRT_LAYER3 = 1'b0; $stop;
    #100;
    $stop;
end

endmodule